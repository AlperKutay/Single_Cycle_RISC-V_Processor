/*
	R-Type: ALU and SHIFT operations
	I-Type: LOAD,SHIFT[I],ALU[I] and JALR operations
	S-Type: STORE opeations
	B-Type: BRANCH operations
	U-Type: LUI and AUIPC operations
	J-Type: JAL operation
*/

module Controller 
	(
		input clk, reset,
		input [31:0]Instr,Zero,
		output reg [3:0]ALUControl, 
		output reg [2:0]ImmSrc,
		output reg PCSrc, ResultSrc, ALUSrc,
		output reg RegWrite, MemWrite,
		output reg [4:0] shamt
	);
	
	localparam	xADD = 4'b0000,
					xSUB = 4'b0001,
					xSLT = 4'b0010,
					xSLTU= 4'b0011,
					xXOR = 4'b0100,
					xORR = 4'b0101,
					xAND = 4'b0110,
					xSLL = 4'b0111,
					xSRL = 4'b1000,
					xSRA = 4'b1001,
					xADDU= 4'b1010,
					xSUBU= 4'b1011;
	
	localparam	ADD_SUB = 3'b000,
					SLL = 3'b001,
					SLT = 3'b010,
					SLTU= 3'b011,
					XOR = 3'b100,
					SRL_SRA = 3'b101,
					ORR = 3'b110,
					AND = 3'b111;
					
	localparam 	ALU_SHIFT = 7'b0110011,
					LOAD = 7'b0000011,
					ALUI_SHIFTI = 7'b0010011,
					JALR = 7'b1100111,
					STORE = 7'b0100011,
					BRANCH = 7'b1100011,
					LUI = 7'b0110111,
					AUIPC = 7'b0010111,
					JAL = 7'b1101111;

	localparam 	R_TYPE = 3'b111,
					I_TYPE = 3'b000,
					S_TYPE = 3'b001,
					B_TYPE = 3'b010,
					U_TYPE = 3'b011,
					J_TYPE = 3'b100;
					
	localparam	LB = 3'b000,
					LH = 3'b001,
					LW = 3'b010,
					LBU= 3'b100,
					LHU= 3'b101;

	localparam	SB = 3'b000,
					SH = 3'b001,
					SW = 3'b010;					
	
	localparam	BEQ = 3'b000,
					BNE = 3'b001,
					BLT = 3'b100,
					BGE = 3'b101,
					BLTU= 3'b110,
					BGEU= 3'b111;
	
	wire [7:0]op;
	wire [2:0]funct3;
	wire funct7_5;
	wire [4:0] rs2,rs1,rd;
	
	assign op = Instr[6:0];
	assign funct3 = Instr[14:12];
	assign funct7_5 = Instr[30];
	assign rs1 = Instr[19:15];
	assign rs2 = Instr[24:20];
	assign rd = Instr[11:7];
	
	always@(*) begin
		
		case(op)
			//R-TYPE
			ALU_SHIFT: begin
				ImmSrc = R_TYPE;
				PCSrc = 1'b0;
				ResultSrc  = 1'b0;
				ALUSrc = 1'b0;
				RegWrite = 1'b1;
				MemWrite = 1'b0;
				shamt = rs2;				
				case(funct3)
					ADD_SUB:begin
						if(funct7_5 == 1'b0) begin //ADD
							ALUControl = xADD;
						end
						else begin						//SUB
							ALUControl = xSUB;					
						end
					end
					SLL:begin						
						ALUControl = xSLL;						
					end
					SLT:begin
						ALUControl = xSLT;					
					end
					SLTU:begin
						ALUControl = xSLTU;					
					end
					XOR:begin
						ALUControl = xXOR;				
					end
					SRL_SRA:begin						
						if(funct7_5 == 1'b0) begin //SRL
							ALUControl = xSRL;							
						end
						else begin						//SRA
							ALUControl = xSRA;							
						end
					end
					ORR:begin				
						ALUControl = xORR;				
					end
					AND:begin					
						ALUControl = xAND;					
					end
				endcase
			end
			//I-TYPE
			LOAD: begin
				ImmSrc = I_TYPE;
				PCSrc = 1'b0;
				ResultSrc  = 1'b1;
				ALUSrc = 1'b1;
				RegWrite = 1'b1;
				MemWrite = 1'b0;
				shamt = rs2;
				case(funct3)
					LB:begin
						ALUControl = xADD;
					end
					LH:begin
						ALUControl = xADD;
					end
					LW:begin
						ALUControl = xADD;
					end
					LBU:begin
						ALUControl = xADDU;
					end
					LHU:begin
						ALUControl = xADDU;
					end
				endcase
			end
			ALUI_SHIFTI: begin
				ImmSrc = I_TYPE;
				PCSrc = 1'b0;
				ResultSrc  = 1'b0;
				ALUSrc = 1'b1;
				RegWrite = 1'b1;
				MemWrite = 1'b0;
				shamt = rs2;				
				case(funct3)
					ADD_SUB:begin
						ALUControl = xADD;			
					end
					SLL:begin						
						ALUControl = xSLL;						
					end
					SLT:begin
						ALUControl = xSLT;					
					end
					SLTU:begin
						ALUControl = xSLTU;					
					end
					XOR:begin
						ALUControl = xXOR;				
					end
					SRL_SRA:begin						
						if(funct7_5 == 1'b0) begin //SRL
							ALUControl = xSRL;							
						end
						else begin						//SRA
							ALUControl = xSRA;							
						end
					end
					ORR:begin				
						ALUControl = xORR;				
					end
					AND:begin					
						ALUControl = xAND;					
					end
				endcase			
			end
		
			JALR: begin
			
			end
			//S-TYPE
			STORE:begin
				ImmSrc = S_TYPE;
				PCSrc = 1'b0;
				ResultSrc  = 1'b0;
				ALUSrc = 1'b1;
				RegWrite = 1'b0;
				MemWrite = 1'b1;
				shamt = rs2;
				case(funct3)
					SB:begin
						ALUControl = xADD;
					end
					SH:begin
						ALUControl = xADD;
					end
					SW:begin
						ALUControl = xADD;
					end
				endcase				
			end
			//B_TYPE
			BRANCH:begin
				ImmSrc = B_TYPE;
				ResultSrc  = 1'b0;
				ALUSrc = 1'b0;
				RegWrite = 1'b0;
				MemWrite = 1'b0;
				shamt = rs2;				
				case(funct3)
					BEQ:begin
						ALUControl = xSUB;
						PCSrc = (Zero == 32'b0)? 1'b1:1'b0;
					end
					BNE:begin
						ALUControl = xSUB;
						PCSrc = (Zero != 32'b0)? 1'b1:1'b0;					
					end
					BLT:begin
						ALUControl = xSUB;
						PCSrc = (Zero < 32'b0)? 1'b1:1'b0;
					end
					BGE:begin
						ALUControl = xSUB;
						PCSrc = (Zero >= 32'b0)? 1'b1:1'b0;
					end
					BLTU:begin
						ALUControl = xSUBU;
						PCSrc = (Zero < 32'b0)? 1'b1:1'b0;
					end
					BGEU:begin
						ALUControl = xSUBU;
						PCSrc = (Zero >= 32'b0)? 1'b1:1'b0;
					end
				endcase
			end
			//U_TYPE
			LUI:begin
			
			end
			
			AUIPC:begin
			
			end
			//J_TYPE
			JAL:begin
			
			end
			
			default: begin
			
			end
		endcase
	end
	
endmodule
